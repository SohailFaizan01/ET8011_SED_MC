Active_E_Field_Probe
C3 2 1 C value={C_s} vinit=0
C4 1 LGref C value={0.5*C_s} vinit=0
M1 LGref 1 0 0 M
M2 LGref 1 0 0 M
R3 LGref out R value=50 noisetemp={T_op_max} noiseflow=0 dcvar=0 dcvarlot=0
R4 out 0 R value=50 noisetemp={T_op_max} noiseflow=0 dcvar=0 dcvarlot=0
V1 2 0 V value={V_in} noise=0 dc=0 dcvar=0
.end