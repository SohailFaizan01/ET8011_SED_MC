Active_E-Field_Probe
C2 4 2 C value={C_s} vinit=0
D1 0 2 D
G1 2 0 1 0 G value=0.5*{C_s}
G2 2 0 3 0 G value=2.5*{C_s}
H1 3 0 5 H value=5
N1 1 3 2 0 N
R2 1 0 R value=50 noisetemp=0 noiseflow=0 dcvar=0 dcvarlot=0
V1 4 0 V value={V_in} noise=0 dc=0 dcvar=0
.end