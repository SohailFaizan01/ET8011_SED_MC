Active_E_Field_Probe
.param V_D=1.8 V_G=0.5 V_S=0 W=10u L=180n
.source V1
.detector V_out
.lgref Gm_M1_X1
C12 1 3 C value={C_s} vinit=0
C13 3 2 C value={0.5*C_s} vinit=0
R6 2 out R value=50 noisetemp={T_op_max} noiseflow=0 dcvar=0 dcvarlot=0
R7 out 0 R value=50 noisetemp={T_op_max} noiseflow=0 dcvar=0 dcvarlot=0
V1 1 0 V value={V_in} noise=0 dc=0 dcvar=0
X1 2 3 0 0 CMOS18N_V W={W} L={L} VG={V_G} VD={V_D} VS={V_S}
.end