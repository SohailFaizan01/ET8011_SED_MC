Active_E_Field_Probe
C1 2 1 C value={C_s} vinit=0
C2 8 Amp_out C value={0.56*C_s} vinit=0
R1 1 8 R value={R_ph} noisetemp={T_op_max} noiseflow=0 dcvar=0 dcvarlot=0
R2 Amp_out vo R value=50 noisetemp={T_op_max} noiseflow=0 dcvar=0 dcvarlot=0
R3 vo 0 R value=50 noisetemp={0} noiseflow=0 dcvar=0 dcvarlot=0
V1 2 0 V value={V_in} noise=0 dc=0 dcvar=0
X1 3 4 5 6 CMOS18ND W={W1_N} L={L1_N} ID={ID1_N}
X2 Amp_out 7 0 0 CMOS18P W={W_P} L={L_P} ID={ID_P}
X3 Amp_out 7 0 0 CMOS18N W={W_N} L={L_N} ID={ID_N}
X4 8 0 5 MN18_noise ID={ID1_N} IG={0} W={W1_N} L={L1_N}
X5 0 0 6 MN18_noise ID={ID1_N} IG={0} W={W1_N} L={L1_N}
X6 0 0 3 0 CMOS18N W={0.025*W1_N} L={L1_N} ID={ID1_N}
X7 7 0 4 0 CMOS18N W={0.025*W1_N} L={L1_N} ID={ID1_N}
.end