Active_E-Field_Probe
C1 3 4 C value=? vinit=0
D1 0 2 D
D2 0 3 D
E1 2 0 1 0 EZ value=? zo=?
N1 1 0 2 0 N
N2 4 0 3 0 N
R1 5 2 R value=? noisetemp=0 noiseflow=0 dcvar=0 dcvarlot=0
R2 0 1 R value=? noisetemp=0 noiseflow=0 dcvar=0 dcvarlot=0
R3 6 3 R value=? noisetemp=0 noiseflow=0 dcvar=0 dcvarlot=0
R4 0 4 R value=? noisetemp=0 noiseflow=0 dcvar=0 dcvarlot=0
V1 5 0 V value=? noise=0 dc=0 dcvar=0
V2 6 0 V value=? noise=0 dc=0 dcvar=0
.end